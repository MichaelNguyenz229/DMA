module dma_desc_fetch
(
    input clk,
    input reset,
)