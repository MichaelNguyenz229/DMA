module dma_write_block
(
    input clk,
    input reset,

    //to AVMM master port
    output [31:0] wr_master_addr_o,
    output [10:0] wr_master_bcount_o,
    output [255:0] wr_master_data_o,

    //from AVMM master port
    input wr_master_wait_req_i,

    //from desc processsor
    input dma_wr_fifo_command_req_i,
    input [15:0] dma_wr_bytes_to_transfer_i,
    input [31:0] dma_wr_addr_i,

    //to desc processor
    output dma_wr_fifo_full_o,

    //to status update block
    output dma_status_fifo_wr_req_o,
    output [24:0] dma_status_fifo_data_o,

    //from status update block
    input dma_status_fifo_almost_full_i,

    //from dma data fifo
    output [255:0] dma_wr_data
);

//internal signals
wire [47:0] wr_fifo_data_in;
wire [47:0] wr_fifo_data_q;

wire wr_fifo_empty;

reg [2:0] current_state;
reg [2:0] next_state;

//write block fifo
scfifo	write_block_fifo (
				.clock (clk),
				.data (wr_fifo_data_in),
				.rdreq (state),
				.sclr (reset),
				.wrreq (dma_wr_fifo_command_req_i),
				.almost_full (),
				.q (wr_fifo_data_q),
				.aclr (),
				.almost_empty (),
				.eccstatus (),
				.empty (wr_fifo_empty),
				.full (dma_wr_fifo_full_o),
				.usedw ());
	defparam
		write_block_fifo.add_ram_output_register = "OFF",
		write_block_fifo.almost_full_value = 24,
		write_block_fifo.intended_device_family = "Cyclone V",
		write_block_fifo.lpm_numwords = 32,
		write_block_fifo.lpm_showahead = "OFF",
		write_block_fifo.lpm_type = "scfifo",
		write_block_fifo.lpm_width = 48,
		write_block_fifo.lpm_widthu = 5,
		write_block_fifo.overflow_checking = "ON",
		write_block_fifo.underflow_checking = "ON",
		write_block_fifo.use_eab = "ON";

//write block state machine
localparam IDLE = 3'b00;
localparam RD_CMD_FIFO = 3'b001;
localparam LD_CMD_REG = 3'b010;
localparam CHECK_XFR = 3'b011;
localparam XFR_DATA = 3'b100;
localparam UPDATE_STATUS = 3'b101;

always @ (posedge clk)
    if(reset)
        current_state <= IDLE;
    else
        current_state <= next_state;

always @*
    case(current_state)
        IDLE:

        RD_CMD_FIFO:

        LD_CMD_REG:

        CHECK_XFR:

        XFR_DATA:

        UPDATE_STATUS:

        default:
        
    endcase

//state machine assignment
assign idle_state = (current_state[2:0] == IDLE);
assign rd_cmd_fifo_state = (current_state[2:0] == RD_CMD_FIFO);
assign ld_cmd_reg_state = (current_state[2:0] == LD_CMD_REG);
assign check_xfr_state = (current_state[2:0] == CHECK_XFR);
assign xfr_data_state = (current_state[2:0] == XFR_DATA);
assign update_status_state = (current_state[2:0] == UPDATE_STATUS);
